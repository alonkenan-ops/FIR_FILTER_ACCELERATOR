`include "defines.svh"

module partial_prod_gen (
    input  logic [15:0] i_sample,
    input  logic [15:0] i_coeff,
    output logic [31:0] o_rows [0:15] // a lot of fucking dots aint it
);

endmodule