`include "defines.svh"

module rounding_sat (
    input  logic [35:0] i_data,
    output logic [15:0] o_data
);

endmodule