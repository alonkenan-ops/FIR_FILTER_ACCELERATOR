`include "defines.svh"

module final_adder (
    input  logic [35:0] i_sum_vec,
    input  logic [35:0] i_carry_vec,
    output logic [35:0] o_result
);

endmodule